
package config_pkg;
    parameter P_DATA_WIDTH = 16,
              P_CLK_DIV    = 4,
              P_CS_POLAR   = 0;
endpackage
