
package config_pkg;
    parameter P_DATA_WIDTH = 8,
              P_CLK_DIV    = 2,
              P_CS_POLAR   = 0;
endpackage
